`timescale 1ns / 1ps

module tb_exponent_comparator;

    

endmodule
