`timescale 1ns / 1ps

module tb_fpu_adder;

    reg clk;
    reg [31:0] a, b;
    reg [1:0] op;
    wire [31:0] out;
    
    fpu_top DUT (.clk(clk),
                 .a(a),
                 .b(b),
                 .op(op),
                 .out(out));
                 
    initial begin
    
        clk = 0;
        op = 2'b00;
        
        //  0.0 + 0.0 = 0.0
        //  out = 0_00000000_00000000000000000000000
        a = 32'b0_00000000_00000000000000000000000;
        b = 32'b0_00000000_00000000000000000000000;
        #50
        
        //  1.25 + 1.50 = 2.75
        //  out = 0_10000000_01100000000000000000000
        //        0_10000101_01100000000000000000000
        a = 32'b0_01111111_01000000000000000000000;
        b = 32'b0_01111111_10000000000000000000000;
        #50
        
        //  43.75 + 5.25 = 49.0
        a = 32'b0_10000100_01011110000000000000000;
        b = 32'b0_10000001_01010000000000000000000;
        #50
    
        $finish;
    end
    
    always #1 clk = ~clk;

endmodule
